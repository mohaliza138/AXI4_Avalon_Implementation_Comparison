module avalon_st_wrapper ();
endmodule
