module axi4_wrapper ();
endmodule
