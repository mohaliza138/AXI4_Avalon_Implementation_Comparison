module avalon_mm_slave_wrapper ();



endmodule
