module axi4_lite_wrapper ();
endmodule
