module axi4_stream_wrapper ();
endmodule
