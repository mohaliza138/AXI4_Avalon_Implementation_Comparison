module avalon_mm_wrapper ();
endmodule
