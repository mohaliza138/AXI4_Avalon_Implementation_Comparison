// `define VERBOSE
